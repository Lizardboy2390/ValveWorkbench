* Triode model

.subckt triode A G1 K
.param MU=112.986
.param KG1=463.667
.param X=1.24465
.param KP=848.497
.param KVB=0.191374
.param KVB1=72.2789
.param VCT=0.361821

R1 G1 K 1G
R2 A K 1G
R3 1 K 1G

EPK 1 K VALUE={pow(V(A,K)*log(1.0+exp(KP*(1.0/MU+(V(G1,K)+VCT)/sqrt(KVB+KVB1*V(A,K)+V(A,K)^2))))/KP,X)}

GA A K VALUE={V(1,K)/KG1}

.ends
