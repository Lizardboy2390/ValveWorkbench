Test harness for biasing pentodes

.include pentode.cir

.param MU=31.9482
.param KG1=998.437
.param X=1.56336
.param KP=167.091
.param KVB=0.000248849
.param KVB1=19.8172
.param VCT=0.0

.param KG2=5655.41
.param A=0.0
.param ALPHA=0.249777
.param BETA=0.0643662
.param GAMMA=0.798651

.param KG2A=6709.55
.param TAU=0.434771
.param RHO=0.0547342
.param THETA=0.854024
.param PSI=4.91385

.param OMEGA=270.473
.param LAMBDA=63.8964
.param NU=29.9968
.param S=0.307751
.param AP=0.00755009

.param OS=-0.000344448

VA 1 0 dc 300
VG2 3 0 dc 140
VM1 1 4 dc 0
VM2 3 5 dc 0

VG1 0 2 dc 0

X1 4 5 2 0 pentode MU={MU} KG1={KG1} X={X} KP={KP} KVB={KVB} KVB1={KVB1} VCT={VCT}
+                  KG2={KG2} A={A} ALPHA={ALPHA} BETA={BETA} GAMMA={GAMMA}
+                  KG2A={KG2A} TAU={TAU} RHO={RHO} THETA={THETA} PSI={PSI}
+                  OMEGA={OMEGA} LAMBDA={LAMBDA} NU={NU} S={S} AP={AP}
+                  OS={OS}

.dc VA 0 300 1 VG1 0 5 0.5

.control

run
plot {I(VM1)} {I(VM2)}

.endc

.end